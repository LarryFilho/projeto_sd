LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

PACKAGE NAO_PACKAGE IS
	COMPONENT NAO
		PORT (x: IN STD_LOGIC_VECTOR(3 DOWNTO 0) ;
					s : OUT STD_LOGIC_VECTOR(3 DOWNTO 0) 
				);
	END COMPONENT;
END NAO_PACKAGE;