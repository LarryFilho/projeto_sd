LIBRARY IEEE ;
USE IEEE.STD_LOGIC_1164.all ;
USE work.FULL_ADDER_PACKAGE.all ;

ENTITY RIPPLE_CARRY IS

	PORT (Cin: IN STD_LOGIC;
				A, B: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
				SAIDA: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
				Cout: OUT STD_LOGIC
			);
				
END RIPPLE_CARRY ;

ARCHITECTURE logica OF RIPPLE_CARRY IS

SIGNAL CARRY_AUXILIAR: STD_LOGIC_VECTOR(3 DOWNTO 0);

SIGNAL AUX: STD_LOGIC_VECTOR(3 DOWNTO 0);


BEGIN

	WITH Cin SELECT
		AUX <= B WHEN '0',
			not B WHEN OTHERS;

	STAGE0: FULLADDER PORT MAP(Cin, 					 A(0), AUX(0), SAIDA(0), CARRY_AUXILIAR(0));
	STAGE1: FULLADDER PORT MAP(CARRY_AUXILIAR(0), A(1), AUX(1), SAIDA(1), CARRY_AUXILIAR(1));
	STAGE2: FULLADDER PORT MAP(CARRY_AUXILIAR(1), A(2), AUX(2), SAIDA(2), CARRY_AUXILIAR(2));
	STAGE3: FULLADDER PORT MAP(CARRY_AUXILIAR(2), A(3), AUX(3), SAIDA(3), Cout);
	
END logica ;