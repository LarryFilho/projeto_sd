LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE work.RIPPLE_CARRY_PACKAGE.all;
USE work.E_PACKAGE.all;
USE work.OU_PACKAGE.all;
USE work.NAO_PACKAGE.all;
USE work.COMPARADOR_PACKAGE.all;

ENTITY ULA IS

	PORT (ALU_OPERATION: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
				A, B: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
				COUT, ZERO, OVERFLOW, EQU, GRT, LST: OUT STD_LOGIC;
				RESULT: OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
			);
				
END ULA ;

ARCHITECTURE logica OF ULA IS

SIGNAL COUT_SOMA, COUT_SUB : STD_LOGIC;

SIGNAL RESULT_SOMA_AUXILIAR: STD_LOGIC_VECTOR(3 DOWNTO 0);

SIGNAL RESULT_SUB_AUXILIAR: STD_LOGIC_VECTOR(3 DOWNTO 0);

SIGNAL RESULT_AND: STD_LOGIC_VECTOR(3 DOWNTO 0);

SIGNAL RESULT_OR: STD_LOGIC_VECTOR(3 DOWNTO 0);

SIGNAL RESULT_NAO: STD_LOGIC_VECTOR(3 DOWNTO 0);

SIGNAL EQU_SIGNAL, GRT_SIGNAL, LST_SIGNAL : STD_LOGIC;

BEGIN

STAGE0: E  PORT MAP(A, B, RESULT_AND);
STAGE1: OU PORT MAP(A, B, RESULT_OR);
STAGE2: NAO PORT MAP(B, RESULT_NAO);
STAGE4: RIPPLE_CARRY PORT MAP('0', A, B, RESULT_SOMA_AUXILIAR, COUT_SOMA);
STAGE5: RIPPLE_CARRY PORT MAP('1', A, B, RESULT_SUB_AUXILIAR, COUT_SUB);
STAGE6: COMPARADOR PORT MAP(A, B, EQU_SIGNAL, GRT_SIGNAL, LST_SIGNAL);

		
RESULT <= "0000" 		WHEN ALU_OPERATION = "000" ELSE
			 RESULT_AND WHEN ALU_OPERATION = "001" ELSE
			 RESULT_OR  WHEN ALU_OPERATION = "010" ELSE
			 RESULT_NAO WHEN ALU_OPERATION = "011" ELSE
			 RESULT_SOMA_AUXILIAR WHEN ALU_OPERATION = "100" ELSE
			 RESULT_SUB_AUXILIAR  WHEN ALU_OPERATION = "101" ELSE
			 (others => 'U');
			 
EQU <= EQU_SIGNAL when ALU_OPERATION = "111" ELSE '0';
GRT <= GRT_SIGNAL when ALU_OPERATION = "111" ELSE '0';
LST <= LST_SIGNAL when ALU_OPERATION = "111" ELSE '0';
	

COUT <= COUT_SOMA WHEN ALU_OPERATION = "100" ELSE			
		  COUT_SUB  WHEN ALU_OPERATION = "101" ELSE 
		  '0';
		  
		  
ZERO <= '1' WHEN (RESULT = "0000" AND ALU_OPERATION /= "000") ELSE '0';


END logica;