LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

PACKAGE OU_PACKAGE IS
	COMPONENT OU
		PORT (x, y : IN STD_LOGIC_VECTOR(3 DOWNTO 0) ;
					s : OUT STD_LOGIC_VECTOR(3 DOWNTO 0) 
				);
	END COMPONENT;
END OU_PACKAGE;