LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

PACKAGE COMPARADOR_PACKAGE IS
	COMPONENT COMPARADOR
		PORT (A, B : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
				EQUAL, GREATER, LESS: OUT STD_LOGIC 
			);
	END COMPONENT;
END COMPARADOR_PACKAGE;