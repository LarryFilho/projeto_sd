LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

PACKAGE ULA_PACKAGE IS
	COMPONENT ULA
		PORT (ALU_OPERATION: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
				A, B: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
				COUT, ZERO, OVERFLOW, EQU, GRT, LST: OUT STD_LOGIC;
				RESULT: OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
			);
	END COMPONENT;
END ULA_PACKAGE;