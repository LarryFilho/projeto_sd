LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

PACKAGE E_PACKAGE IS
	COMPONENT E
		PORT (x, y : IN STD_LOGIC_VECTOR(3 DOWNTO 0) ;
				s : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
				);
	END COMPONENT;
END E_PACKAGE;