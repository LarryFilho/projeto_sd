LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL ;
USE IEEE.STD_LOGIC_SIGNED.ALL;

ENTITY E IS
	
	PORT (x, y : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
				s : OUT STD_LOGIC_VECTOR(3 DOWNTO 0) 
			);
	END E ;

ARCHITECTURE logica OF E IS

BEGIN

	s <= x AND y;


END logica ;