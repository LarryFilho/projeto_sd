LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL ;
USE IEEE.STD_LOGIC_SIGNED.ALL;

ENTITY NAO IS
	
	PORT (x: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
				s : OUT STD_LOGIC_VECTOR(3 DOWNTO 0) 
			);
	END NAO ;

ARCHITECTURE logica OF NAO IS

BEGIN

	s <= NOT X;


END logica ;