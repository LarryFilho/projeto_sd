LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

PACKAGE FULL_ADDER_PACKAGE IS
	COMPONENT FULLADDER
		PORT(Cin, x, y: in STD_LOGIC;
				s, Cout : OUT STD_LOGIC
			 );
	END COMPONENT;
END FULL_ADDER_PACKAGE;