LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

PACKAGE RIPPLE_CARRY_PACKAGE IS
	COMPONENT RIPPLE_CARRY
		PORT (Cin: IN STD_LOGIC;
				A, B: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
				SAIDA: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
				Cout: OUT STD_LOGIC
			);
	END COMPONENT;
END RIPPLE_CARRY_PACKAGE;